LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY Exercicio_3 IS
	PORT (	A: IN std_logic_vector(1 downto 0);
	     SAIDA: OUT std_logic_vector(1 downto 0));
END Exercicio_3;

ARCHITECTURE logica OF Exercicio_3 IS
	SIGNAL 

BEGIN
	SAIDA : 
END logica;