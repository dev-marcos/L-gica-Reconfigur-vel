LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY Exercicio_1 IS
	PORT (	A: IN std_logic_vector(1 downto 0);
	     SAIDA: OUT std_logic_vector(1 downto 0));
END Exercicio_1;

ARCHITECTURE logica OF Exercicio_1 IS
	SIGNAL 

BEGIN
	SAIDA : 
END logica;