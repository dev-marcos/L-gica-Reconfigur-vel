LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY Exercicio_2 IS
	PORT (	A: IN std_logic_vector(1 downto 0);
	     SAIDA: OUT std_logic_vector(1 downto 0));
END Exercicio_2;

ARCHITECTURE logica OF Exercicio_2 IS
	SIGNAL 

BEGIN
	SAIDA : 
END logica;