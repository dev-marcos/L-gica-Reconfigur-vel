LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY Exercicio_4 IS
	PORT (	 A: IN std_logic;
				 B: IN std_logic; 
				EN: IN std_logic;
			  SUM: OUT std_logic;
			 COUT: OUT std_logic;

END Exercicio_4;

ARCHITECTURE logica OF Exercicio_4 IS
SIGNAL 

BEGIN
	SUM : 
	
	
END logica;